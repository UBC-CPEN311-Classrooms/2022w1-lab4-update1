module tb_rtl_wordcopy();
endmodule: tb_rtl_wordcopy
