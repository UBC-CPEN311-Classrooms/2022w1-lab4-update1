module tb_rtl_dot();
endmodule: tb_rtl_dot
