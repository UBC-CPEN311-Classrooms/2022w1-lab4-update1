module tb_vga_avalon();

// Your testbench goes here.

endmodule: tb_vga_avalon
